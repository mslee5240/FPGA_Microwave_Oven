`timescale 1ns / 1ps

//==============================================================================
// 클럭 분주기 모듈 - 100MHz를 1Hz로 분주
// 동작 원리: 카운터 기반 토글 방식으로 정확한 1초 주기 클럭 생성
// 용도: 전자레인지 타이머의 1초 단위 카운트다운용
//==============================================================================
module clock_divider(
    input clk,              // 100MHz 시스템 클럭 (BASYS-3 보드 기본 클럭)
    input reset,            // 비동기 리셋 (Active High)
    output reg clk_1hz      // 1Hz 출력 클럭 (1초마다 토글)
);

    //==========================================================================
    // 분주 비율 계산
    // 100MHz → 1Hz: 100,000,000:1 분주 필요
    // 토글 방식: 반주기(0.5초)마다 토글하여 1초 주기 생성
    // 따라서 50,000,000 카운트마다 토글 = 1Hz 클럭 생성
    //==========================================================================
    parameter COUNT_MAX = 50_000_000 - 1;      // 49,999,999까지 카운트
    
    // 50,000,000을 카운트하기 위한 카운터
    // 2^26 = 67,108,864 > 50,000,000 이므로 26비트면 충분
    reg [25:0] counter = 0;
    
    //==========================================================================
    // 메인 분주 로직 - 100MHz 클럭에 동기화
    //==========================================================================
    always @(posedge clk, posedge reset) begin
        if (reset) begin
            // 리셋 시 초기화: 카운터와 출력 클럭을 0으로 설정
            counter <= 0;
            clk_1hz <= 0;
        end else begin
            // 50,000,000 카운트 완료 시 (정확히 0.5초 경과)
            if (counter == COUNT_MAX) begin
                counter <= 0;              // 카운터 리셋
                clk_1hz <= ~clk_1hz;       // 출력 클럭 토글 (0→1 또는 1→0)
            end else begin
                // 아직 0.5초가 안 됨: 카운터 계속 증가
                counter <= counter + 1;
            end
        end
    end

    //==========================================================================
    // 동작 타이밍 설명:
    // - 매 클럭(10ns)마다 카운터 +1
    // - 49,999,999까지 카운트 = 500,000,000ns = 0.5초
    // - 0.5초마다 clk_1hz 토글 = 1초 주기 완성
    // - 결과: 듀티 사이클 50%의 정확한 1Hz 클럭 출력
    //==========================================================================

endmodule